// Verilog netlist created by Tang Dynasty v5.6.71036
// Mon Oct  2 10:49:58 2023

`timescale 1ns / 1ps
module atan
  (
  clk,
  rst,
  start,
  xin,
  yin,
  angle,
  done
  );

  input clk;
  input rst;
  input start;
  input [17:0] xin;
  input [17:0] yin;
  output [18:0] angle;
  output done;

  parameter COMPENSATION = "No Compensation";
  parameter ITERATION = 16;
  parameter PRECISION = 16;
  parameter SCALED = 0;
  // localparam PI = 19'b0110010010000111111;
  // localparam W_CNT = 5;
  wire [18:0] al_63c792c7;
  wire [18:0] al_67a58a3a;
  wire [19:0] al_a9c1cf7a;
  wire [19:0] al_fa21b72a;
  wire [19:0] al_86bba01f;
  wire [19:0] al_d670b90a;
  wire [4:0] al_a3e2b42;
  wire [4:0] al_55146f8b;
  wire [4:0] al_b029b709;
  wire [4:0] al_2ca2eaaa;
  wire [16:0] al_43ee5b62;
  wire [16:0] al_a8a039bd;
  wire [17:0] al_655add9;
  wire [17:0] al_bb54b22f;
  wire [17:0] al_aa605bd8;
  wire [17:0] al_e8eb449b;
  wire [17:0] al_8145a529;
  wire [17:0] al_f178cf22;
  wire [17:0] al_ba2f1510;
  wire [17:0] al_615e209b;
  wire [17:0] al_e890342d;
  wire [17:0] al_b0aa8206;
  wire [17:0] al_f774eaf9;
  wire [17:0] al_8b1ee5d9;
  wire [17:0] al_12c226aa;
  wire [17:0] al_7b6549fa;
  wire [17:0] al_54f6e7c3;
  wire [17:0] al_d6af4c70;
  wire [17:0] al_a89eb1ca;
  wire [17:0] al_deeec3ed;
  wire [17:0] al_9a3f7017;
  wire [17:0] al_9addee19;
  wire al_2d23a90d;
  wire al_a6a3e0a0;
  wire al_1140b89f;
  wire al_aa18e7c5;
  wire al_b4e29609;
  wire al_4c46f7ea;
  wire al_2c776044;
  wire al_912aa5d5;
  wire al_49b15ec;
  wire al_d05c69c9;
  wire al_64d14f69;
  wire al_312b3af4;
  wire al_1f0013fa;
  wire al_99f44ac;
  wire al_d0045161;
  wire al_16c52ec8;
  wire al_af21225a;
  wire al_8ba9d093;
  wire al_d2041f17;
  wire al_477219c8;
  wire al_df76032a;
  wire al_ff46c763;
  wire al_a22e7e39;
  wire al_54d446b6;
  wire al_6e13aef1;
  wire al_afc156cf;
  wire al_c0326560;
  wire al_eb56e8c8;
  wire al_c703b21a;
  wire al_f2295687;
  wire al_ea857007;
  wire al_a3d28a21;
  wire al_8edb520a;
  wire al_103cd50f;
  wire al_8b138a0b;
  wire al_b322bc2;
  wire al_c483235b;
  wire al_cbb4d2e8;
  wire al_f48b56af;
  wire al_a651a3d3;
  wire al_50aa345c;
  wire al_bad9c600;
  wire al_3f2ceda0;
  wire al_2b36ec4c;
  wire al_beaff734;
  wire al_11f09a69;
  wire al_90e32614;
  wire al_771e9c44;
  wire al_64588870;
  wire al_86e106a8;
  wire al_25036e36;
  wire al_e99edde6;
  wire al_bb47cbad;
  wire al_4a06208;
  wire al_1eb004f0;
  wire al_f96e4e54;
  wire al_10d96161;
  wire al_f62f8727;
  wire al_ca754152;
  wire al_8a2de5e1;
  wire al_1e6d359a;
  wire al_7cb51e63;
  wire al_88ae6f58;
  wire al_7de19a8c;
  wire al_e75e71a9;
  wire al_60eb3689;
  wire al_f6fb6313;
  wire al_6cce137;
  wire al_db44397d;
  wire al_f3df5f83;
  wire al_cdcf1edb;
  wire al_2788f29f;
  wire al_9ce8bde4;
  wire al_3b7e2483;
  wire al_f66288b;
  wire al_ee2cc5d5;
  wire al_6b105db6;
  wire al_e2334515;
  wire al_b25ed4d7;
  wire al_a8c455aa;
  wire al_6fffff50;
  wire al_7dc82f77;
  wire al_e8c1ab1e;
  wire al_1af2bab3;
  wire al_60dcbcf6;
  wire al_f4e90bd7;
  wire al_d4f4ffd4;
  wire al_4c0923e5;
  wire al_794e2cf3;
  wire al_3c6b7670;
  wire al_ad05e543;
  wire al_397f5efc;
  wire al_64bfb744;
  wire al_c5a5deba;
  wire al_661904d9;
  wire al_be443a52;
  wire al_6d594c9b;
  wire al_2c6ea385;
  wire al_ce6e5997;
  wire al_1f65ec13;
  wire al_11fe6cd4;
  wire al_40b705d7;
  wire al_a743530c;
  wire al_a5be61f4;
  wire al_f577d7c;
  wire al_f39a7e9;
  wire al_9762a925;
  wire al_ef2ad0c3;
  wire al_e7f7dbb1;
  wire al_b1f223c3;
  wire al_e7086bfe;
  wire al_5e7e4908;
  wire al_d16993ed;
  wire al_ae0a6293;
  wire al_d07a623a;
  wire al_126bbf82;
  wire al_1aac3445;
  wire al_f5516224;
  wire al_91108e0e;
  wire al_a4e1781b;
  wire al_dc44be48;
  wire al_d8dd00e3;
  wire al_a0bad8f5;
  wire al_daf1c16d;
  wire al_24d9d8b6;
  wire al_4ff4ec95;
  wire al_e54de9c;
  wire al_583f8393;
  wire al_4d59c3c7;
  wire al_216911ff;
  wire al_93ee307b;
  wire al_c1faafeb;
  wire al_c6d867e6;
  wire al_1041605;
  wire al_b59343a1;
  wire al_fb401a7e;
  wire al_54e68679;
  wire al_bbe72ea1;
  wire al_ae3b43d5;
  wire al_9d2e2c47;
  wire al_a525c35;
  wire al_99de34c9;
  wire al_1271c79c;
  wire al_a129eed6;
  wire al_81880b1d;
  wire al_14e87bc7;
  wire al_51ec8425;
  wire al_2bd93fd7;
  wire al_7830f36d;
  wire al_254eb4e8;
  wire al_deb4d477;
  wire al_4d3cc22;
  wire al_916512e5;
  wire al_d5f320f0;
  wire al_8b75dfd4;
  wire al_67ea5570;
  wire al_54208fc4;
  wire al_99cfa891;
  wire al_31bcf06d;
  wire al_cd305354;
  wire al_5f6ba172;
  wire al_83a98034;
  wire al_543f4953;
  wire al_c6d22991;
  wire al_c04f33dd;
  wire al_3379f791;
  wire al_803879c7;
  wire al_48cbf9af;
  wire al_4f9f19b;
  wire al_5a076585;
  wire al_1ce14aac;
  wire al_854c573f;
  wire al_c03651db;
  wire al_73eda6f6;
  wire al_747e69b3;
  wire al_51f316f6;
  wire al_8a394456;
  wire al_9047c71;
  wire al_1259ba86;
  wire al_9800fd32;
  wire al_af16dfa7;
  wire al_87b4efd6;
  wire al_1f3b4767;
  wire al_4ab15cc0;
  wire al_86baf6c6;
  wire al_abf6101b;
  wire al_a26df073;
  wire al_75f92221;
  wire al_60b812b4;
  wire al_b5005b7;
  wire al_895351d0;
  wire al_e841d7a8;
  wire al_e08923c5;
  wire al_45f63f66;
  wire al_5072ec3a;
  wire al_64522de4;
  wire al_6bd097c8;
  wire al_489ab129;
  wire al_d32b8d83;
  wire al_e54f5937;
  wire al_267693c3;
  wire al_f2ea1b91;
  wire al_185cfc7b;
  wire al_ab37028c;
  wire al_c41ea483;
  wire al_40edf471;
  wire al_14d0775;
  wire al_e0531380;
  wire al_3c344131;
  wire al_88f2b0ea;
  wire al_923aa1f3;
  wire al_4c309c76;
  wire al_2b296468;
  wire al_9ea7dc42;
  wire al_e7e648ec;
  wire al_c18c443d;
  wire al_879333c8;
  wire al_63f07c7f;
  wire al_f120ad54;
  wire al_72ad6500;
  wire al_b2a8a0cc;
  wire al_80739918;
  wire al_67d43207;
  wire al_f42f533c;
  wire al_853b0020;
  wire al_6c78c52c;
  wire al_598dbbb7;
  wire al_a2275c94;
  wire al_1fb8f7d6;
  wire al_137b074e;
  wire al_6d3f1d3d;
  wire al_2013c010;
  wire al_22d6ddd;
  wire al_b5596380;
  wire al_65737be6;
  wire al_967be913;
  wire al_dce5c03c;
  wire al_48b19352;
  wire al_fb209166;
  wire al_b77cbcd0;
  wire al_6075e6a9;
  wire al_492fb484;
  wire al_248f265c;
  wire al_efe81361;
  wire al_1de057dc;
  wire al_399025e4;
  wire al_6652589d;
  wire al_9aa2c63b;
  wire al_44f78eb0;
  wire al_b494668c;
  wire al_96795d02;
  wire al_85347eda;
  wire al_2853bf2a;
  wire al_ce27e68f;
  wire al_5f96adf7;
  wire al_c29dd627;
  wire al_31cf9bca;
  wire al_329701d8;
  wire al_9ca1c07c;
  wire al_d92048f7;
  wire al_6af624ab;
  wire al_4772cc8e;
  wire al_1883443;
  wire al_dee61509;
  wire al_ce078ee;
  wire al_2b0d498c;

  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c22ee456 (
    .a(al_a9c1cf7a[5]),
    .b(al_43ee5b62[5]),
    .c(al_912aa5d5),
    .o({al_49b15ec,al_86bba01f[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4f8c6b2 (
    .a(al_a9c1cf7a[6]),
    .b(al_43ee5b62[6]),
    .c(al_49b15ec),
    .o({al_d05c69c9,al_86bba01f[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_251c9501 (
    .a(al_a9c1cf7a[7]),
    .b(al_43ee5b62[7]),
    .c(al_d05c69c9),
    .o({al_64d14f69,al_86bba01f[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b10f851 (
    .a(al_a9c1cf7a[8]),
    .b(al_43ee5b62[8]),
    .c(al_64d14f69),
    .o({al_312b3af4,al_86bba01f[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f6074d25 (
    .a(al_a9c1cf7a[9]),
    .b(al_43ee5b62[9]),
    .c(al_312b3af4),
    .o({al_1f0013fa,al_86bba01f[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_fa8db078 (
    .a(al_a9c1cf7a[10]),
    .b(al_43ee5b62[10]),
    .c(al_1f0013fa),
    .o({al_99f44ac,al_86bba01f[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_77855a53 (
    .a(al_a9c1cf7a[11]),
    .b(al_43ee5b62[11]),
    .c(al_99f44ac),
    .o({al_d0045161,al_86bba01f[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e3fa0367 (
    .a(al_a9c1cf7a[12]),
    .b(al_43ee5b62[12]),
    .c(al_d0045161),
    .o({al_16c52ec8,al_86bba01f[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f953a96c (
    .a(al_a9c1cf7a[13]),
    .b(al_43ee5b62[13]),
    .c(al_16c52ec8),
    .o({al_af21225a,al_86bba01f[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_65c8a090 (
    .a(al_a9c1cf7a[14]),
    .b(al_43ee5b62[14]),
    .c(al_af21225a),
    .o({al_8ba9d093,al_86bba01f[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_53b7c044 (
    .a(al_a9c1cf7a[15]),
    .b(al_43ee5b62[15]),
    .c(al_8ba9d093),
    .o({al_d2041f17,al_86bba01f[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d4fabdf4 (
    .a(al_a9c1cf7a[16]),
    .b(1'b0),
    .c(al_d2041f17),
    .o({al_477219c8,al_86bba01f[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4c333d3d (
    .a(al_a9c1cf7a[17]),
    .b(1'b0),
    .c(al_477219c8),
    .o({al_df76032a,al_86bba01f[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ad500350 (
    .a(al_a9c1cf7a[18]),
    .b(1'b0),
    .c(al_df76032a),
    .o({al_ff46c763,al_86bba01f[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d576b9a4 (
    .a(al_a9c1cf7a[19]),
    .b(1'b0),
    .c(al_ff46c763),
    .o({open_n0,al_86bba01f[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_cda14380 (
    .a(1'b0),
    .o({al_1140b89f,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f54c3dbb (
    .a(al_a9c1cf7a[0]),
    .b(al_43ee5b62[0]),
    .c(al_1140b89f),
    .o({al_aa18e7c5,al_86bba01f[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c9b145c3 (
    .a(al_a9c1cf7a[1]),
    .b(al_43ee5b62[1]),
    .c(al_aa18e7c5),
    .o({al_b4e29609,al_86bba01f[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_85743617 (
    .a(al_a9c1cf7a[2]),
    .b(al_43ee5b62[2]),
    .c(al_b4e29609),
    .o({al_4c46f7ea,al_86bba01f[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ad670f93 (
    .a(al_a9c1cf7a[3]),
    .b(al_43ee5b62[3]),
    .c(al_4c46f7ea),
    .o({al_2c776044,al_86bba01f[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ec16458c (
    .a(al_a9c1cf7a[4]),
    .b(al_43ee5b62[4]),
    .c(al_2c776044),
    .o({al_912aa5d5,al_86bba01f[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_2165f23d (
    .a(1'b0),
    .o({al_a22e7e39,open_n6}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_5a77c71d (
    .a(al_f178cf22[8]),
    .b(al_9addee19[8]),
    .c(al_ea857007),
    .o({al_a3d28a21,al_615e209b[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_6113318c (
    .a(al_f178cf22[9]),
    .b(al_9addee19[9]),
    .c(al_a3d28a21),
    .o({al_8edb520a,al_615e209b[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1ba0daa2 (
    .a(al_f178cf22[10]),
    .b(al_9addee19[10]),
    .c(al_8edb520a),
    .o({al_103cd50f,al_615e209b[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4ff26d7e (
    .a(al_f178cf22[11]),
    .b(al_9addee19[11]),
    .c(al_103cd50f),
    .o({al_8b138a0b,al_615e209b[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b257243f (
    .a(al_f178cf22[12]),
    .b(al_9addee19[12]),
    .c(al_8b138a0b),
    .o({al_b322bc2,al_615e209b[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_ce1cc971 (
    .a(al_f178cf22[13]),
    .b(al_9addee19[13]),
    .c(al_b322bc2),
    .o({al_c483235b,al_615e209b[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e3dc02b8 (
    .a(al_f178cf22[14]),
    .b(al_9addee19[14]),
    .c(al_c483235b),
    .o({al_cbb4d2e8,al_615e209b[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9fa2507d (
    .a(al_f178cf22[15]),
    .b(al_9addee19[15]),
    .c(al_cbb4d2e8),
    .o({al_f48b56af,al_615e209b[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f7236576 (
    .a(al_f178cf22[16]),
    .b(al_9addee19[16]),
    .c(al_f48b56af),
    .o({al_a651a3d3,al_615e209b[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_d5b75486 (
    .a(al_f178cf22[17]),
    .b(al_d6af4c70[17]),
    .c(al_a651a3d3),
    .o({open_n7,al_615e209b[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_61c46b5d (
    .a(al_f178cf22[0]),
    .b(al_9addee19[0]),
    .c(al_a22e7e39),
    .o({al_54d446b6,al_615e209b[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9c5c9996 (
    .a(al_f178cf22[1]),
    .b(al_9addee19[1]),
    .c(al_54d446b6),
    .o({al_6e13aef1,al_615e209b[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c04cf982 (
    .a(al_f178cf22[2]),
    .b(al_9addee19[2]),
    .c(al_6e13aef1),
    .o({al_afc156cf,al_615e209b[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f1d55d58 (
    .a(al_f178cf22[3]),
    .b(al_9addee19[3]),
    .c(al_afc156cf),
    .o({al_c0326560,al_615e209b[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_212b0a99 (
    .a(al_f178cf22[4]),
    .b(al_9addee19[4]),
    .c(al_c0326560),
    .o({al_eb56e8c8,al_615e209b[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_4a0be642 (
    .a(al_f178cf22[5]),
    .b(al_9addee19[5]),
    .c(al_eb56e8c8),
    .o({al_c703b21a,al_615e209b[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_9d22fee2 (
    .a(al_f178cf22[6]),
    .b(al_9addee19[6]),
    .c(al_c703b21a),
    .o({al_f2295687,al_615e209b[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a9fc3313 (
    .a(al_f178cf22[7]),
    .b(al_9addee19[7]),
    .c(al_f2295687),
    .o({al_ea857007,al_615e209b[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    al_6c65e6ec (
    .a(1'b0),
    .o({al_50aa345c,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7a814cc1 (
    .a(al_d6af4c70[8]),
    .b(al_b0aa8206[8]),
    .c(al_64588870),
    .o({al_86e106a8,al_9a3f7017[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_3f0f1414 (
    .a(al_d6af4c70[9]),
    .b(al_b0aa8206[9]),
    .c(al_86e106a8),
    .o({al_25036e36,al_9a3f7017[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_bd625e74 (
    .a(al_d6af4c70[10]),
    .b(al_b0aa8206[10]),
    .c(al_25036e36),
    .o({al_e99edde6,al_9a3f7017[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f66cc420 (
    .a(al_d6af4c70[11]),
    .b(al_b0aa8206[11]),
    .c(al_e99edde6),
    .o({al_bb47cbad,al_9a3f7017[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_be113f82 (
    .a(al_d6af4c70[12]),
    .b(al_b0aa8206[12]),
    .c(al_bb47cbad),
    .o({al_4a06208,al_9a3f7017[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_197ca113 (
    .a(al_d6af4c70[13]),
    .b(al_b0aa8206[13]),
    .c(al_4a06208),
    .o({al_1eb004f0,al_9a3f7017[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_16c07b12 (
    .a(al_d6af4c70[14]),
    .b(al_b0aa8206[14]),
    .c(al_1eb004f0),
    .o({al_f96e4e54,al_9a3f7017[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_e77d29a3 (
    .a(al_d6af4c70[15]),
    .b(al_b0aa8206[15]),
    .c(al_f96e4e54),
    .o({al_10d96161,al_9a3f7017[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_a710bda1 (
    .a(al_d6af4c70[16]),
    .b(al_b0aa8206[16]),
    .c(al_10d96161),
    .o({al_f62f8727,al_9a3f7017[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_21783b3a (
    .a(al_d6af4c70[17]),
    .b(al_f178cf22[17]),
    .c(al_f62f8727),
    .o({open_n11,al_9a3f7017[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c2cd2d4e (
    .a(al_d6af4c70[0]),
    .b(al_b0aa8206[0]),
    .c(al_50aa345c),
    .o({al_bad9c600,al_9a3f7017[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_39375266 (
    .a(al_d6af4c70[1]),
    .b(al_b0aa8206[1]),
    .c(al_bad9c600),
    .o({al_3f2ceda0,al_9a3f7017[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_1be482f2 (
    .a(al_d6af4c70[2]),
    .b(al_b0aa8206[2]),
    .c(al_3f2ceda0),
    .o({al_2b36ec4c,al_9a3f7017[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_63d33a4b (
    .a(al_d6af4c70[3]),
    .b(al_b0aa8206[3]),
    .c(al_2b36ec4c),
    .o({al_beaff734,al_9a3f7017[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_c797f8a4 (
    .a(al_d6af4c70[4]),
    .b(al_b0aa8206[4]),
    .c(al_beaff734),
    .o({al_11f09a69,al_9a3f7017[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_7f656e5 (
    .a(al_d6af4c70[5]),
    .b(al_b0aa8206[5]),
    .c(al_11f09a69),
    .o({al_90e32614,al_9a3f7017[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_b11b3677 (
    .a(al_d6af4c70[6]),
    .b(al_b0aa8206[6]),
    .c(al_90e32614),
    .o({al_771e9c44,al_9a3f7017[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    al_f1a11535 (
    .a(al_d6af4c70[7]),
    .b(al_b0aa8206[7]),
    .c(al_771e9c44),
    .o({al_64588870,al_9a3f7017[7]}));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_74f9489f (
    .a(al_86bba01f[0]),
    .b(al_67a58a3a[0]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[0]),
    .o(al_fa21b72a[0]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_fa1c403b (
    .a(al_86bba01f[10]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[10]),
    .o(al_fa21b72a[10]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_bca178ce (
    .a(al_86bba01f[11]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[11]),
    .o(al_fa21b72a[11]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_3f45dbda (
    .a(al_86bba01f[12]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[12]),
    .o(al_fa21b72a[12]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_e4ef7c04 (
    .a(al_86bba01f[13]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[13]),
    .o(al_fa21b72a[13]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_c5ad99f (
    .a(al_86bba01f[14]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[14]),
    .o(al_fa21b72a[14]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_b58571f9 (
    .a(al_86bba01f[15]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[15]),
    .o(al_fa21b72a[15]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_45d470a2 (
    .a(al_86bba01f[16]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[16]),
    .o(al_fa21b72a[16]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_b24c5c3b (
    .a(al_86bba01f[17]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[17]),
    .o(al_fa21b72a[17]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_b21fd745 (
    .a(al_86bba01f[18]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[18]),
    .o(al_fa21b72a[18]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_2a973b65 (
    .a(al_86bba01f[19]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[19]),
    .o(al_fa21b72a[19]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_5ef4cb6 (
    .a(al_86bba01f[1]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[1]),
    .o(al_fa21b72a[1]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_11e2dce1 (
    .a(al_86bba01f[2]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[2]),
    .o(al_fa21b72a[2]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_6455bad3 (
    .a(al_86bba01f[3]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[3]),
    .o(al_fa21b72a[3]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_90ed3722 (
    .a(al_86bba01f[4]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[4]),
    .o(al_fa21b72a[4]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_eabd8aaf (
    .a(al_86bba01f[5]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[5]),
    .o(al_fa21b72a[5]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_acf00b84 (
    .a(al_86bba01f[6]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[6]),
    .o(al_fa21b72a[6]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_4fa713e1 (
    .a(al_86bba01f[7]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[7]),
    .o(al_fa21b72a[7]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_1af0e313 (
    .a(al_86bba01f[8]),
    .b(al_67a58a3a[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[8]),
    .o(al_fa21b72a[8]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'hccfacc0a))
    al_dfd46c01 (
    .a(al_86bba01f[9]),
    .b(al_67a58a3a[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_d670b90a[9]),
    .o(al_fa21b72a[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_1c1ac75 (
    .a(al_5a076585),
    .b(al_1ce14aac),
    .c(al_b029b709[4]),
    .o(al_543f4953));
  AL_DFF_X al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_543f4953),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_7583f4d6 (
    .a(al_b029b709[3]),
    .b(al_b029b709[4]),
    .o(al_cd305354));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_3765d349 (
    .a(al_b029b709[1]),
    .b(al_b029b709[2]),
    .o(al_c04f33dd));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~(~C*~(B*A))))"),
    .INIT(32'h00ff0007))
    al_a5f59856 (
    .a(al_cd305354),
    .b(al_c04f33dd),
    .c(al_b029b709[0]),
    .d(al_48cbf9af),
    .e(al_4f9f19b),
    .o(al_2ca2eaaa[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*(B@A))"),
    .INIT(16'h0006))
    al_566b91ed (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_48cbf9af),
    .d(al_4f9f19b),
    .o(al_2ca2eaaa[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*(C@(B*A)))"),
    .INIT(32'h00000078))
    al_b6c49bd1 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_48cbf9af),
    .e(al_4f9f19b),
    .o(al_2ca2eaaa[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*B*A))"),
    .INIT(16'h807f))
    al_d573f520 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_c6d22991));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_5caaf660 (
    .a(al_c6d22991),
    .b(al_48cbf9af),
    .c(al_4f9f19b),
    .o(al_2ca2eaaa[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_2b9b0b78 (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_a6a3e0a0));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*(B@A))"),
    .INIT(16'h0006))
    al_ca573301 (
    .a(al_a6a3e0a0),
    .b(al_b029b709[4]),
    .c(al_48cbf9af),
    .d(al_4f9f19b),
    .o(al_2ca2eaaa[4]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_1f11638d (
    .a(al_a8a039bd[14]),
    .b(al_a3e2b42[0]),
    .o(al_ca754152));
  AL_MAP_LUT5 #(
    .EQN("(~A*~B*~C*~D*~E+A*~B*~C*~D*~E+A*B*~C*~D*~E+A*~B*C*~D*~E+~A*B*C*~D*~E+A*B*C*~D*~E+~A*~B*~C*D*~E+A*~B*~C*D*~E+~A*B*~C*D*~E+A*B*~C*D*~E+~A*~B*C*D*~E+A*~B*C*D*~E+~A*B*C*D*~E+A*B*C*D*~E+~A*~B*~C*~D*E)"),
    .INIT(32'b00000000000000011111111111101011))
    al_38df2f87 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .e(al_a3e2b42[4]),
    .o(al_a8a039bd[0]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_83686079 (
    .a(1'b0),
    .o({al_8a2de5e1,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5dce2a87 (
    .a(1'b0),
    .b(yin[8]),
    .c(al_6cce137),
    .o({al_db44397d,al_aa605bd8[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6016763 (
    .a(1'b0),
    .b(yin[9]),
    .c(al_db44397d),
    .o({al_f3df5f83,al_aa605bd8[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d632c6d (
    .a(1'b0),
    .b(yin[10]),
    .c(al_f3df5f83),
    .o({al_cdcf1edb,al_aa605bd8[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b4fa7b84 (
    .a(1'b0),
    .b(yin[11]),
    .c(al_cdcf1edb),
    .o({al_2788f29f,al_aa605bd8[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_76976ed5 (
    .a(1'b0),
    .b(yin[12]),
    .c(al_2788f29f),
    .o({al_9ce8bde4,al_aa605bd8[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acf7562e (
    .a(1'b0),
    .b(yin[13]),
    .c(al_9ce8bde4),
    .o({al_3b7e2483,al_aa605bd8[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e853baae (
    .a(1'b0),
    .b(yin[14]),
    .c(al_3b7e2483),
    .o({al_f66288b,al_aa605bd8[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72dfb0ec (
    .a(1'b0),
    .b(yin[15]),
    .c(al_f66288b),
    .o({al_ee2cc5d5,al_aa605bd8[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d348c1c8 (
    .a(1'b0),
    .b(yin[16]),
    .c(al_ee2cc5d5),
    .o({al_6b105db6,al_aa605bd8[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f294e788 (
    .a(1'b0),
    .b(yin[17]),
    .c(al_6b105db6),
    .o({open_n15,al_aa605bd8[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b24fb310 (
    .a(1'b0),
    .b(yin[0]),
    .c(al_8a2de5e1),
    .o({al_1e6d359a,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f7bda68 (
    .a(1'b0),
    .b(yin[1]),
    .c(al_1e6d359a),
    .o({al_7cb51e63,al_aa605bd8[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e0f5d561 (
    .a(1'b0),
    .b(yin[2]),
    .c(al_7cb51e63),
    .o({al_88ae6f58,al_aa605bd8[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be99a96b (
    .a(1'b0),
    .b(yin[3]),
    .c(al_88ae6f58),
    .o({al_7de19a8c,al_aa605bd8[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2bd3c09b (
    .a(1'b0),
    .b(yin[4]),
    .c(al_7de19a8c),
    .o({al_e75e71a9,al_aa605bd8[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_65a5e647 (
    .a(1'b0),
    .b(yin[5]),
    .c(al_e75e71a9),
    .o({al_60eb3689,al_aa605bd8[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff6ca422 (
    .a(1'b0),
    .b(yin[6]),
    .c(al_60eb3689),
    .o({al_f6fb6313,al_aa605bd8[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d02400f (
    .a(1'b0),
    .b(yin[7]),
    .c(al_f6fb6313),
    .o({al_6cce137,al_aa605bd8[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_fb918c26 (
    .a(1'b0),
    .o({al_e2334515,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5c76d5bb (
    .a(1'b0),
    .b(al_655add9[8]),
    .c(al_f4e90bd7),
    .o({al_d4f4ffd4,al_54f6e7c3[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c052b85 (
    .a(1'b0),
    .b(al_655add9[9]),
    .c(al_d4f4ffd4),
    .o({al_4c0923e5,al_54f6e7c3[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_44b78d1 (
    .a(1'b0),
    .b(al_655add9[10]),
    .c(al_4c0923e5),
    .o({al_794e2cf3,al_54f6e7c3[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_99955157 (
    .a(1'b0),
    .b(al_655add9[11]),
    .c(al_794e2cf3),
    .o({al_3c6b7670,al_54f6e7c3[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8170adb (
    .a(1'b0),
    .b(al_655add9[12]),
    .c(al_3c6b7670),
    .o({al_ad05e543,al_54f6e7c3[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54f5eb45 (
    .a(1'b0),
    .b(al_655add9[13]),
    .c(al_ad05e543),
    .o({al_397f5efc,al_54f6e7c3[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41596a54 (
    .a(1'b0),
    .b(al_655add9[14]),
    .c(al_397f5efc),
    .o({al_64bfb744,al_54f6e7c3[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_19439718 (
    .a(1'b0),
    .b(al_655add9[15]),
    .c(al_64bfb744),
    .o({al_c5a5deba,al_54f6e7c3[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd6e9ba (
    .a(1'b0),
    .b(al_655add9[16]),
    .c(al_c5a5deba),
    .o({al_661904d9,al_54f6e7c3[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37173e61 (
    .a(1'b0),
    .b(al_655add9[17]),
    .c(al_661904d9),
    .o({open_n20,al_54f6e7c3[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_afe79d12 (
    .a(1'b0),
    .b(al_655add9[0]),
    .c(al_e2334515),
    .o({al_b25ed4d7,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2823027 (
    .a(1'b0),
    .b(al_655add9[1]),
    .c(al_b25ed4d7),
    .o({al_a8c455aa,al_54f6e7c3[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ab4ef237 (
    .a(1'b0),
    .b(al_655add9[2]),
    .c(al_a8c455aa),
    .o({al_6fffff50,al_54f6e7c3[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73b14a62 (
    .a(1'b0),
    .b(al_655add9[3]),
    .c(al_6fffff50),
    .o({al_7dc82f77,al_54f6e7c3[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59c31ac2 (
    .a(1'b0),
    .b(al_655add9[4]),
    .c(al_7dc82f77),
    .o({al_e8c1ab1e,al_54f6e7c3[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae30f0a9 (
    .a(1'b0),
    .b(al_655add9[5]),
    .c(al_e8c1ab1e),
    .o({al_1af2bab3,al_54f6e7c3[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f518f82 (
    .a(1'b0),
    .b(al_655add9[6]),
    .c(al_1af2bab3),
    .o({al_60dcbcf6,al_54f6e7c3[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fce5a731 (
    .a(1'b0),
    .b(al_655add9[7]),
    .c(al_60dcbcf6),
    .o({al_f4e90bd7,al_54f6e7c3[7]}));
  AL_DFF_X al_e2342da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5f6ba172),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_63c792c7[8]));
  AL_DFF_X al_795dec5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[8]));
  AL_DFF_X al_e8b27f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[9]));
  AL_DFF_X al_34c43e91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[10]));
  AL_DFF_X al_4034d121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[11]));
  AL_DFF_X al_7260e525 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[12]));
  AL_DFF_X al_c152e5cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[13]));
  AL_DFF_X al_6e95db6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[14]));
  AL_DFF_X al_58944ff2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[15]));
  AL_DFF_X al_22fef235 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[16]));
  AL_DFF_X al_7d508833 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(yin[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[17]));
  AL_DFF_X al_6eb318e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[0]));
  AL_DFF_X al_10074c95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[1]));
  AL_DFF_X al_5fb1cf51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[2]));
  AL_DFF_X al_dc5daab3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[3]));
  AL_DFF_X al_5394044a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[4]));
  AL_DFF_X al_b89d9b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[5]));
  AL_DFF_X al_81c5ed9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[6]));
  AL_DFF_X al_9e15c642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b1ee5d9[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f774eaf9[7]));
  AL_DFF_X al_c26c9bb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[8]));
  AL_DFF_X al_7256805c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[9]));
  AL_DFF_X al_3579341e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[10]));
  AL_DFF_X al_b7079f11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[11]));
  AL_DFF_X al_89cb7fac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[12]));
  AL_DFF_X al_7f48cb2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[13]));
  AL_DFF_X al_8c60f702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[14]));
  AL_DFF_X al_2e772330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[15]));
  AL_DFF_X al_835d154d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[16]));
  AL_DFF_X al_d32f36bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[17]));
  AL_DFF_X al_de040350 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[0]));
  AL_DFF_X al_25378cfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[1]));
  AL_DFF_X al_dc93576e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[2]));
  AL_DFF_X al_76b20766 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[3]));
  AL_DFF_X al_a8ce422 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[4]));
  AL_DFF_X al_e3895fe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[5]));
  AL_DFF_X al_2160ccea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[6]));
  AL_DFF_X al_df8e007c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7b6549fa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_12c226aa[7]));
  AL_DFF_X al_b40a42c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[8]));
  AL_DFF_X al_56fbb473 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[9]));
  AL_DFF_X al_f912cfa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[10]));
  AL_DFF_X al_790357b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[11]));
  AL_DFF_X al_1f745e25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[12]));
  AL_DFF_X al_fdf3d1b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[13]));
  AL_DFF_X al_28c56aa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[14]));
  AL_DFF_X al_fa1f6a4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[15]));
  AL_DFF_X al_7852efc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[16]));
  AL_DFF_X al_9a72719d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[17]));
  AL_DFF_X al_31c2c18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[0]));
  AL_DFF_X al_bed75354 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[1]));
  AL_DFF_X al_b2c2a4b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[2]));
  AL_DFF_X al_99383aba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[3]));
  AL_DFF_X al_f8178b2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[4]));
  AL_DFF_X al_be1fc3e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[5]));
  AL_DFF_X al_c9f8b2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[6]));
  AL_DFF_X al_5979435b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a89eb1ca[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6af4c70[7]));
  AL_DFF_X al_b40e8e05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be443a52),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67a58a3a[8]));
  AL_DFF_X al_2259e8d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a98034),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67a58a3a[9]));
  AL_DFF_X al_fd544ba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6d594c9b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67a58a3a[0]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    al_5e95843a (
    .a(al_83a98034),
    .b(al_63c792c7[8]),
    .o(al_6d594c9b));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_d701a9b8 (
    .a(al_83a98034),
    .b(al_63c792c7[8]),
    .o(al_be443a52));
  AL_DFF_X al_596b0fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[8]));
  AL_DFF_X al_5cfa2c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[9]));
  AL_DFF_X al_c56c02f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[10]));
  AL_DFF_X al_60ec2662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[11]));
  AL_DFF_X al_ea3f598e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[12]));
  AL_DFF_X al_dd4ae85d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[13]));
  AL_DFF_X al_e2aa8055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[14]));
  AL_DFF_X al_82aa8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[15]));
  AL_DFF_X al_7f911c70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[16]));
  AL_DFF_X al_8908ba38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[17]));
  AL_DFF_X al_16ad90bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[0]));
  AL_DFF_X al_2149b062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[18]));
  AL_DFF_X al_56d82898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[19]));
  AL_DFF_X al_e1044ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[1]));
  AL_DFF_X al_16da6de4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[2]));
  AL_DFF_X al_e819e904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[3]));
  AL_DFF_X al_4990808d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[4]));
  AL_DFF_X al_d51e17ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[5]));
  AL_DFF_X al_b67f884b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[6]));
  AL_DFF_X al_ff3308ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fa21b72a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a9c1cf7a[7]));
  AL_DFF_X al_c1e3ea45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[8]));
  AL_DFF_X al_b7aa029f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[9]));
  AL_DFF_X al_2f4f18cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[10]));
  AL_DFF_X al_42a7eb97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[11]));
  AL_DFF_X al_f77c099a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[12]));
  AL_DFF_X al_6893ba8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[13]));
  AL_DFF_X al_d6d1e991 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[14]));
  AL_DFF_X al_4d3bf6cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[15]));
  AL_DFF_X al_aa8c310 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[16]));
  AL_DFF_X al_d8095998 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[17]));
  AL_DFF_X al_53efe64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[0]));
  AL_DFF_X al_68082bd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[18]));
  AL_DFF_X al_26890f76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[1]));
  AL_DFF_X al_802c7023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[2]));
  AL_DFF_X al_9c45670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[3]));
  AL_DFF_X al_b0a0e999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[4]));
  AL_DFF_X al_739d9f2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[5]));
  AL_DFF_X al_7f9eee7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[6]));
  AL_DFF_X al_741313a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9c1cf7a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(angle[7]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_cbb21b57 (
    .a(al_a3e2b42[3]),
    .b(al_a3e2b42[4]),
    .o(al_a743530c));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_50032887 (
    .a(al_a743530c),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .o(al_a8a039bd[14]));
  AL_DFF_X al_5e904a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_40b705d7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3e2b42[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*(B@A))"),
    .INIT(16'h0006))
    al_db3b2b53 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_803879c7),
    .d(al_48cbf9af),
    .o(al_2c6ea385));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*(C@(B*A)))"),
    .INIT(32'h00000078))
    al_4496adb2 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_803879c7),
    .e(al_48cbf9af),
    .o(al_ce6e5997));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_db38e2c4 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .o(al_2d23a90d));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*A))"),
    .INIT(16'h7f80))
    al_b910420c (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .o(al_55146f8b[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_90d7e42b (
    .a(al_55146f8b[3]),
    .b(al_803879c7),
    .c(al_48cbf9af),
    .o(al_1f65ec13));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*(B@A))"),
    .INIT(16'h0006))
    al_f16a60a9 (
    .a(al_2d23a90d),
    .b(al_a3e2b42[4]),
    .c(al_803879c7),
    .d(al_48cbf9af),
    .o(al_11fe6cd4));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~D*~(~B*~A)))"),
    .INIT(16'h0f01))
    al_91adf23 (
    .a(al_a8a039bd[14]),
    .b(al_a3e2b42[0]),
    .c(al_803879c7),
    .d(al_48cbf9af),
    .o(al_40b705d7));
  AL_DFF_X al_116f1db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c6ea385),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3e2b42[1]));
  AL_DFF_X al_6c993e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce6e5997),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3e2b42[2]));
  AL_DFF_X al_23963ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1f65ec13),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3e2b42[3]));
  AL_DFF_X al_6c25cf29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_11fe6cd4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a3e2b42[4]));
  AL_DFF_X al_cbbb4490 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2ca2eaaa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[0]));
  AL_DFF_X al_30153836 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2ca2eaaa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[1]));
  AL_DFF_X al_37ead40d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2ca2eaaa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[2]));
  AL_DFF_X al_7625712c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2ca2eaaa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[3]));
  AL_DFF_X al_2531de5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_2ca2eaaa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b029b709[4]));
  AL_DFF_X al_3b229c23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[8]));
  AL_DFF_X al_cf6e7591 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[9]));
  AL_DFF_X al_5a2f8048 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[10]));
  AL_DFF_X al_1abb3ac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[11]));
  AL_DFF_X al_78a4a9ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[12]));
  AL_DFF_X al_65b6d202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[13]));
  AL_DFF_X al_647eb39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[14]));
  AL_DFF_X al_369b90e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ca754152),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[15]));
  AL_DFF_X al_139c5590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[0]));
  AL_DFF_X al_39f4cfe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[1]));
  AL_DFF_X al_164ed6d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[2]));
  AL_DFF_X al_2d1248a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[3]));
  AL_DFF_X al_d8e1e88b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[4]));
  AL_DFF_X al_f380c478 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[5]));
  AL_DFF_X al_22301a07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[6]));
  AL_DFF_X al_b389eb27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a8a039bd[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_43ee5b62[7]));
  AL_DFF_X al_db0079e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[8]));
  AL_DFF_X al_876f7db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[9]));
  AL_DFF_X al_69a0ebce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[10]));
  AL_DFF_X al_a6c89e95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[11]));
  AL_DFF_X al_f3acd144 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[12]));
  AL_DFF_X al_f6a3bd12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[13]));
  AL_DFF_X al_22c71420 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[14]));
  AL_DFF_X al_32b9df1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[15]));
  AL_DFF_X al_93449db5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[16]));
  AL_DFF_X al_4ad3d5d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[17]));
  AL_DFF_X al_e87e6f9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[0]));
  AL_DFF_X al_43ae41e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[1]));
  AL_DFF_X al_32098dc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[2]));
  AL_DFF_X al_1771790f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[3]));
  AL_DFF_X al_4e0fd4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[4]));
  AL_DFF_X al_1d1fe749 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[5]));
  AL_DFF_X al_f8b279ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[6]));
  AL_DFF_X al_75a93bc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bb54b22f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_655add9[7]));
  AL_DFF_X al_8117d99a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[8]));
  AL_DFF_X al_170fafe0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[9]));
  AL_DFF_X al_d7229bc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[10]));
  AL_DFF_X al_d80ca115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[11]));
  AL_DFF_X al_a73edca8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[12]));
  AL_DFF_X al_e38dfe07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[13]));
  AL_DFF_X al_3e2268e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[14]));
  AL_DFF_X al_9bbe1751 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[15]));
  AL_DFF_X al_71f8ee87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[16]));
  AL_DFF_X al_619c7086 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[17]));
  AL_DFF_X al_2e8a2570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[0]));
  AL_DFF_X al_4c05617e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[1]));
  AL_DFF_X al_7cbb1b5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[2]));
  AL_DFF_X al_1851373 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[3]));
  AL_DFF_X al_6ef4721c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[4]));
  AL_DFF_X al_ef14836c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[5]));
  AL_DFF_X al_29111b42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[6]));
  AL_DFF_X al_9e5c600b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8145a529[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e8eb449b[7]));
  AL_DFF_X al_8ff57d60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[8]));
  AL_DFF_X al_47b511ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[9]));
  AL_DFF_X al_89005d1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[10]));
  AL_DFF_X al_f5b5ca38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[11]));
  AL_DFF_X al_7907a48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[12]));
  AL_DFF_X al_f3e31ce5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[13]));
  AL_DFF_X al_55389588 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[14]));
  AL_DFF_X al_dc2b1ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[15]));
  AL_DFF_X al_220615c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[16]));
  AL_DFF_X al_c7aa6b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[17]));
  AL_DFF_X al_3176eb22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[0]));
  AL_DFF_X al_1ec04f80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[1]));
  AL_DFF_X al_ec2280f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[2]));
  AL_DFF_X al_ecb5afd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[3]));
  AL_DFF_X al_d15fb662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[4]));
  AL_DFF_X al_e22992ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[5]));
  AL_DFF_X al_c3bb0c4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[6]));
  AL_DFF_X al_5b797485 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ba2f1510[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f178cf22[7]));
  AL_DFF_X al_dce734fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(start),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_803879c7));
  AL_DFF_X al_d5515080 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_803879c7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_48cbf9af));
  AL_DFF_X al_d59b3527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_48cbf9af),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4f9f19b));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b9c8457 (
    .a(al_a9c1cf7a[5]),
    .b(al_43ee5b62[5]),
    .c(al_e7f7dbb1),
    .o({al_b1f223c3,al_d670b90a[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e613dd7 (
    .a(al_a9c1cf7a[6]),
    .b(al_43ee5b62[6]),
    .c(al_b1f223c3),
    .o({al_e7086bfe,al_d670b90a[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27c8842d (
    .a(al_a9c1cf7a[7]),
    .b(al_43ee5b62[7]),
    .c(al_e7086bfe),
    .o({al_5e7e4908,al_d670b90a[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_462a01f1 (
    .a(al_a9c1cf7a[8]),
    .b(al_43ee5b62[8]),
    .c(al_5e7e4908),
    .o({al_d16993ed,al_d670b90a[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b3bce39 (
    .a(al_a9c1cf7a[9]),
    .b(al_43ee5b62[9]),
    .c(al_d16993ed),
    .o({al_ae0a6293,al_d670b90a[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f829bb24 (
    .a(al_a9c1cf7a[10]),
    .b(al_43ee5b62[10]),
    .c(al_ae0a6293),
    .o({al_d07a623a,al_d670b90a[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc29264d (
    .a(al_a9c1cf7a[11]),
    .b(al_43ee5b62[11]),
    .c(al_d07a623a),
    .o({al_126bbf82,al_d670b90a[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee4a1d93 (
    .a(al_a9c1cf7a[12]),
    .b(al_43ee5b62[12]),
    .c(al_126bbf82),
    .o({al_1aac3445,al_d670b90a[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_154312aa (
    .a(al_a9c1cf7a[13]),
    .b(al_43ee5b62[13]),
    .c(al_1aac3445),
    .o({al_f5516224,al_d670b90a[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17566e78 (
    .a(al_a9c1cf7a[14]),
    .b(al_43ee5b62[14]),
    .c(al_f5516224),
    .o({al_91108e0e,al_d670b90a[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_38657e34 (
    .a(al_a9c1cf7a[15]),
    .b(al_43ee5b62[15]),
    .c(al_91108e0e),
    .o({al_a4e1781b,al_d670b90a[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bbcbdbe (
    .a(al_a9c1cf7a[16]),
    .b(1'b0),
    .c(al_a4e1781b),
    .o({al_dc44be48,al_d670b90a[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_216ec453 (
    .a(al_a9c1cf7a[17]),
    .b(1'b0),
    .c(al_dc44be48),
    .o({al_d8dd00e3,al_d670b90a[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c943a4d2 (
    .a(al_a9c1cf7a[18]),
    .b(1'b0),
    .c(al_d8dd00e3),
    .o({al_a0bad8f5,al_d670b90a[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_920ee641 (
    .a(al_a9c1cf7a[19]),
    .b(1'b0),
    .c(al_a0bad8f5),
    .o({open_n22,al_d670b90a[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_68abff86 (
    .a(1'b0),
    .o({al_a5be61f4,open_n25}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8de058bd (
    .a(al_a9c1cf7a[0]),
    .b(al_43ee5b62[0]),
    .c(al_a5be61f4),
    .o({al_f577d7c,al_d670b90a[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbd4c846 (
    .a(al_a9c1cf7a[1]),
    .b(al_43ee5b62[1]),
    .c(al_f577d7c),
    .o({al_f39a7e9,al_d670b90a[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222b6767 (
    .a(al_a9c1cf7a[2]),
    .b(al_43ee5b62[2]),
    .c(al_f39a7e9),
    .o({al_9762a925,al_d670b90a[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c7fbfa5 (
    .a(al_a9c1cf7a[3]),
    .b(al_43ee5b62[3]),
    .c(al_9762a925),
    .o({al_ef2ad0c3,al_d670b90a[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd218d47 (
    .a(al_a9c1cf7a[4]),
    .b(al_43ee5b62[4]),
    .c(al_ef2ad0c3),
    .o({al_e7f7dbb1,al_d670b90a[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_3a3a68e0 (
    .a(1'b0),
    .o({al_daf1c16d,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7a9fe52 (
    .a(al_f178cf22[8]),
    .b(al_9addee19[8]),
    .c(al_c1faafeb),
    .o({al_c6d867e6,al_e890342d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5542edfe (
    .a(al_f178cf22[9]),
    .b(al_9addee19[9]),
    .c(al_c6d867e6),
    .o({al_1041605,al_e890342d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_488602ff (
    .a(al_f178cf22[10]),
    .b(al_9addee19[10]),
    .c(al_1041605),
    .o({al_b59343a1,al_e890342d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5e1d0a51 (
    .a(al_f178cf22[11]),
    .b(al_9addee19[11]),
    .c(al_b59343a1),
    .o({al_fb401a7e,al_e890342d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a28406e8 (
    .a(al_f178cf22[12]),
    .b(al_9addee19[12]),
    .c(al_fb401a7e),
    .o({al_54e68679,al_e890342d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6b74b0b2 (
    .a(al_f178cf22[13]),
    .b(al_9addee19[13]),
    .c(al_54e68679),
    .o({al_bbe72ea1,al_e890342d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_225d9869 (
    .a(al_f178cf22[14]),
    .b(al_9addee19[14]),
    .c(al_bbe72ea1),
    .o({al_ae3b43d5,al_e890342d[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57140763 (
    .a(al_f178cf22[15]),
    .b(al_9addee19[15]),
    .c(al_ae3b43d5),
    .o({al_9d2e2c47,al_e890342d[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2faa1616 (
    .a(al_f178cf22[16]),
    .b(al_9addee19[16]),
    .c(al_9d2e2c47),
    .o({al_a525c35,al_e890342d[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed62317d (
    .a(al_f178cf22[17]),
    .b(al_d6af4c70[17]),
    .c(al_a525c35),
    .o({open_n29,al_e890342d[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5194f578 (
    .a(al_f178cf22[0]),
    .b(al_9addee19[0]),
    .c(al_daf1c16d),
    .o({al_24d9d8b6,al_e890342d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5250c82 (
    .a(al_f178cf22[1]),
    .b(al_9addee19[1]),
    .c(al_24d9d8b6),
    .o({al_4ff4ec95,al_e890342d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce5b7c47 (
    .a(al_f178cf22[2]),
    .b(al_9addee19[2]),
    .c(al_4ff4ec95),
    .o({al_e54de9c,al_e890342d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2348e63f (
    .a(al_f178cf22[3]),
    .b(al_9addee19[3]),
    .c(al_e54de9c),
    .o({al_583f8393,al_e890342d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1dde6515 (
    .a(al_f178cf22[4]),
    .b(al_9addee19[4]),
    .c(al_583f8393),
    .o({al_4d59c3c7,al_e890342d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_730170d3 (
    .a(al_f178cf22[5]),
    .b(al_9addee19[5]),
    .c(al_4d59c3c7),
    .o({al_216911ff,al_e890342d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_81729e9d (
    .a(al_f178cf22[6]),
    .b(al_9addee19[6]),
    .c(al_216911ff),
    .o({al_93ee307b,al_e890342d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73503454 (
    .a(al_f178cf22[7]),
    .b(al_9addee19[7]),
    .c(al_93ee307b),
    .o({al_c1faafeb,al_e890342d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_69abf9ec (
    .a(1'b0),
    .o({al_99de34c9,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dfdc771 (
    .a(al_d6af4c70[8]),
    .b(al_b0aa8206[8]),
    .c(al_254eb4e8),
    .o({al_deb4d477,al_deeec3ed[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e93dcd8b (
    .a(al_d6af4c70[9]),
    .b(al_b0aa8206[9]),
    .c(al_deb4d477),
    .o({al_4d3cc22,al_deeec3ed[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f94769 (
    .a(al_d6af4c70[10]),
    .b(al_b0aa8206[10]),
    .c(al_4d3cc22),
    .o({al_916512e5,al_deeec3ed[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18f640ef (
    .a(al_d6af4c70[11]),
    .b(al_b0aa8206[11]),
    .c(al_916512e5),
    .o({al_d5f320f0,al_deeec3ed[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86ec8670 (
    .a(al_d6af4c70[12]),
    .b(al_b0aa8206[12]),
    .c(al_d5f320f0),
    .o({al_8b75dfd4,al_deeec3ed[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6df03772 (
    .a(al_d6af4c70[13]),
    .b(al_b0aa8206[13]),
    .c(al_8b75dfd4),
    .o({al_67ea5570,al_deeec3ed[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45f02cda (
    .a(al_d6af4c70[14]),
    .b(al_b0aa8206[14]),
    .c(al_67ea5570),
    .o({al_54208fc4,al_deeec3ed[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6b2c7c5 (
    .a(al_d6af4c70[15]),
    .b(al_b0aa8206[15]),
    .c(al_54208fc4),
    .o({al_99cfa891,al_deeec3ed[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86f06d29 (
    .a(al_d6af4c70[16]),
    .b(al_b0aa8206[16]),
    .c(al_99cfa891),
    .o({al_31bcf06d,al_deeec3ed[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff64c9f9 (
    .a(al_d6af4c70[17]),
    .b(al_f178cf22[17]),
    .c(al_31bcf06d),
    .o({open_n33,al_deeec3ed[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6219435f (
    .a(al_d6af4c70[0]),
    .b(al_b0aa8206[0]),
    .c(al_99de34c9),
    .o({al_1271c79c,al_deeec3ed[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9173b3c2 (
    .a(al_d6af4c70[1]),
    .b(al_b0aa8206[1]),
    .c(al_1271c79c),
    .o({al_a129eed6,al_deeec3ed[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e14f1c1 (
    .a(al_d6af4c70[2]),
    .b(al_b0aa8206[2]),
    .c(al_a129eed6),
    .o({al_81880b1d,al_deeec3ed[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b174dbc (
    .a(al_d6af4c70[3]),
    .b(al_b0aa8206[3]),
    .c(al_81880b1d),
    .o({al_14e87bc7,al_deeec3ed[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6657a45b (
    .a(al_d6af4c70[4]),
    .b(al_b0aa8206[4]),
    .c(al_14e87bc7),
    .o({al_51ec8425,al_deeec3ed[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17e08140 (
    .a(al_d6af4c70[5]),
    .b(al_b0aa8206[5]),
    .c(al_51ec8425),
    .o({al_2bd93fd7,al_deeec3ed[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e94e10ff (
    .a(al_d6af4c70[6]),
    .b(al_b0aa8206[6]),
    .c(al_2bd93fd7),
    .o({al_7830f36d,al_deeec3ed[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_440a3abe (
    .a(al_d6af4c70[7]),
    .b(al_b0aa8206[7]),
    .c(al_7830f36d),
    .o({al_254eb4e8,al_deeec3ed[7]}));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+~(B)*~(C)*D+B*~(C)*D))"),
    .INIT(16'h0aa8))
    al_e4ae0e93 (
    .a(al_a743530c),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .d(al_a3e2b42[2]),
    .o(al_a8a039bd[10]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .INIT(16'h02a2))
    al_cc235f61 (
    .a(al_a743530c),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .d(al_a3e2b42[2]),
    .o(al_a8a039bd[11]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_dc1fe16 (
    .a(al_a743530c),
    .b(al_3379f791),
    .c(al_a3e2b42[2]),
    .o(al_a8a039bd[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    al_5a16a101 (
    .a(al_a8a039bd[12]),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .o(al_a8a039bd[13]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*(~(B)*~(C)*~(D)+B*~(C)*~(D)+B*C*D)))"),
    .INIT(32'h00007ff5))
    al_12cf90d1 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .e(al_a3e2b42[4]),
    .o(al_a8a039bd[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D))"),
    .INIT(32'h00003fed))
    al_ac639d52 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .e(al_a3e2b42[4]),
    .o(al_a8a039bd[2]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C@B)))"),
    .INIT(16'h00be))
    al_2ec69993 (
    .a(al_3379f791),
    .b(al_a3e2b42[2]),
    .c(al_a3e2b42[3]),
    .d(al_a3e2b42[4]),
    .o(al_a8a039bd[3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    al_ac52bf53 (
    .a(al_a8a039bd[4]),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .d(al_a3e2b42[2]),
    .o(al_a8a039bd[5]));
  AL_MAP_LUT5 #(
    .EQN("(~E*(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D))"),
    .INIT(32'h000003f8))
    al_74b08c9a (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .c(al_a3e2b42[2]),
    .d(al_a3e2b42[3]),
    .e(al_a3e2b42[4]),
    .o(al_a8a039bd[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_f48539f9 (
    .a(al_a3e2b42[0]),
    .b(al_a3e2b42[1]),
    .o(al_3379f791));
  AL_MAP_LUT4 #(
    .EQN("(~D*(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C))"),
    .INIT(16'h003d))
    al_bd6a53b6 (
    .a(al_3379f791),
    .b(al_a3e2b42[2]),
    .c(al_a3e2b42[3]),
    .d(al_a3e2b42[4]),
    .o(al_a8a039bd[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    al_cc102ffc (
    .a(al_a8a039bd[4]),
    .b(al_a743530c),
    .c(al_3379f791),
    .o(al_a8a039bd[7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*(C@B)))"),
    .INIT(16'haa82))
    al_595cbdf6 (
    .a(al_a743530c),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .d(al_a3e2b42[2]),
    .o(al_a8a039bd[8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(B*~(C)*~(D)+~(B)*C*~(D)+B*C*~(D)+~(B)*~(C)*D+B*~(C)*D+~(B)*C*D))"),
    .INIT(16'h2aa8))
    al_d310e3ed (
    .a(al_a743530c),
    .b(al_a3e2b42[0]),
    .c(al_a3e2b42[1]),
    .d(al_a3e2b42[2]),
    .o(al_a8a039bd[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9953730 (
    .a(al_5f6ba172),
    .b(xin[0]),
    .c(yin[0]),
    .o(al_bb54b22f[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b1cc8be2 (
    .a(al_5f6ba172),
    .b(xin[10]),
    .c(al_aa605bd8[10]),
    .o(al_bb54b22f[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_23b89a4f (
    .a(al_5f6ba172),
    .b(xin[11]),
    .c(al_aa605bd8[11]),
    .o(al_bb54b22f[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e2cb0af1 (
    .a(al_5f6ba172),
    .b(xin[12]),
    .c(al_aa605bd8[12]),
    .o(al_bb54b22f[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fb5002a5 (
    .a(al_5f6ba172),
    .b(xin[13]),
    .c(al_aa605bd8[13]),
    .o(al_bb54b22f[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f80f41af (
    .a(al_5f6ba172),
    .b(xin[14]),
    .c(al_aa605bd8[14]),
    .o(al_bb54b22f[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_80f41a2f (
    .a(al_5f6ba172),
    .b(xin[15]),
    .c(al_aa605bd8[15]),
    .o(al_bb54b22f[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_db9b3c58 (
    .a(al_5f6ba172),
    .b(xin[16]),
    .c(al_aa605bd8[16]),
    .o(al_bb54b22f[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    al_a7dae1c3 (
    .a(xin[17]),
    .b(yin[17]),
    .c(al_aa605bd8[17]),
    .o(al_bb54b22f[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f029d9 (
    .a(al_5f6ba172),
    .b(xin[1]),
    .c(al_aa605bd8[1]),
    .o(al_bb54b22f[1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5263b937 (
    .a(al_5f6ba172),
    .b(xin[2]),
    .c(al_aa605bd8[2]),
    .o(al_bb54b22f[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8c02f654 (
    .a(al_5f6ba172),
    .b(xin[3]),
    .c(al_aa605bd8[3]),
    .o(al_bb54b22f[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1b72b08f (
    .a(al_5f6ba172),
    .b(xin[4]),
    .c(al_aa605bd8[4]),
    .o(al_bb54b22f[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_78d2b06f (
    .a(al_5f6ba172),
    .b(xin[5]),
    .c(al_aa605bd8[5]),
    .o(al_bb54b22f[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d9aee132 (
    .a(al_5f6ba172),
    .b(xin[6]),
    .c(al_aa605bd8[6]),
    .o(al_bb54b22f[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ac3c0d9c (
    .a(al_5f6ba172),
    .b(xin[7]),
    .c(al_aa605bd8[7]),
    .o(al_bb54b22f[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad6d4275 (
    .a(al_5f6ba172),
    .b(xin[8]),
    .c(al_aa605bd8[8]),
    .o(al_bb54b22f[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_286b6fb7 (
    .a(al_5f6ba172),
    .b(xin[9]),
    .c(al_aa605bd8[9]),
    .o(al_bb54b22f[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1357a5a6 (
    .a(al_83a98034),
    .b(al_f774eaf9[0]),
    .c(al_655add9[0]),
    .o(al_8145a529[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_445e91b2 (
    .a(al_83a98034),
    .b(al_f774eaf9[10]),
    .c(al_655add9[10]),
    .o(al_8145a529[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e3b0019a (
    .a(al_83a98034),
    .b(al_f774eaf9[11]),
    .c(al_655add9[11]),
    .o(al_8145a529[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fadf54c5 (
    .a(al_83a98034),
    .b(al_f774eaf9[12]),
    .c(al_655add9[12]),
    .o(al_8145a529[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bc881c1d (
    .a(al_83a98034),
    .b(al_f774eaf9[13]),
    .c(al_655add9[13]),
    .o(al_8145a529[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_e7e7db5b (
    .a(al_83a98034),
    .b(al_f774eaf9[14]),
    .c(al_655add9[14]),
    .o(al_8145a529[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bfce09fc (
    .a(al_83a98034),
    .b(al_f774eaf9[15]),
    .c(al_655add9[15]),
    .o(al_8145a529[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_372e2bc6 (
    .a(al_f774eaf9[17]),
    .b(al_655add9[17]),
    .o(al_83a98034));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c79f5885 (
    .a(al_83a98034),
    .b(al_f774eaf9[16]),
    .c(al_655add9[16]),
    .o(al_8145a529[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_86e1c42c (
    .a(al_f774eaf9[17]),
    .b(al_655add9[17]),
    .o(al_8145a529[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_93acbe72 (
    .a(al_83a98034),
    .b(al_f774eaf9[1]),
    .c(al_655add9[1]),
    .o(al_8145a529[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2333a53b (
    .a(al_83a98034),
    .b(al_f774eaf9[2]),
    .c(al_655add9[2]),
    .o(al_8145a529[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2898e8fd (
    .a(al_83a98034),
    .b(al_f774eaf9[3]),
    .c(al_655add9[3]),
    .o(al_8145a529[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6b6426cc (
    .a(al_83a98034),
    .b(al_f774eaf9[4]),
    .c(al_655add9[4]),
    .o(al_8145a529[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d6d66190 (
    .a(al_83a98034),
    .b(al_f774eaf9[5]),
    .c(al_655add9[5]),
    .o(al_8145a529[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_80b82fe1 (
    .a(al_83a98034),
    .b(al_f774eaf9[6]),
    .c(al_655add9[6]),
    .o(al_8145a529[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a225564b (
    .a(al_83a98034),
    .b(al_f774eaf9[7]),
    .c(al_655add9[7]),
    .o(al_8145a529[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fc0e777d (
    .a(al_83a98034),
    .b(al_f774eaf9[8]),
    .c(al_655add9[8]),
    .o(al_8145a529[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_86fa6982 (
    .a(al_83a98034),
    .b(al_f774eaf9[9]),
    .c(al_655add9[9]),
    .o(al_8145a529[9]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_45ce10c0 (
    .a(al_615e209b[0]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[0]),
    .d(al_48cbf9af),
    .e(al_e890342d[0]),
    .o(al_ba2f1510[0]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_b6c1d5cd (
    .a(al_615e209b[10]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[10]),
    .d(al_48cbf9af),
    .e(al_e890342d[10]),
    .o(al_ba2f1510[10]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_a69939ed (
    .a(al_615e209b[11]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[11]),
    .d(al_48cbf9af),
    .e(al_e890342d[11]),
    .o(al_ba2f1510[11]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_2209fcd7 (
    .a(al_615e209b[12]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[12]),
    .d(al_48cbf9af),
    .e(al_e890342d[12]),
    .o(al_ba2f1510[12]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_9b22f65c (
    .a(al_615e209b[13]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[13]),
    .d(al_48cbf9af),
    .e(al_e890342d[13]),
    .o(al_ba2f1510[13]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_92a221f3 (
    .a(al_615e209b[14]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[14]),
    .d(al_48cbf9af),
    .e(al_e890342d[14]),
    .o(al_ba2f1510[14]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_deab9ae4 (
    .a(al_615e209b[15]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[15]),
    .d(al_48cbf9af),
    .e(al_e890342d[15]),
    .o(al_ba2f1510[15]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_b00a9eff (
    .a(al_615e209b[16]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[16]),
    .d(al_48cbf9af),
    .e(al_e890342d[16]),
    .o(al_ba2f1510[16]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_7f833953 (
    .a(al_615e209b[17]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[17]),
    .d(al_48cbf9af),
    .e(al_e890342d[17]),
    .o(al_ba2f1510[17]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_74a6ddea (
    .a(al_615e209b[1]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[1]),
    .d(al_48cbf9af),
    .e(al_e890342d[1]),
    .o(al_ba2f1510[1]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_4feebaf9 (
    .a(al_615e209b[2]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[2]),
    .d(al_48cbf9af),
    .e(al_e890342d[2]),
    .o(al_ba2f1510[2]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_b41119aa (
    .a(al_615e209b[3]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[3]),
    .d(al_48cbf9af),
    .e(al_e890342d[3]),
    .o(al_ba2f1510[3]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_aae42909 (
    .a(al_615e209b[4]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[4]),
    .d(al_48cbf9af),
    .e(al_e890342d[4]),
    .o(al_ba2f1510[4]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_ef0e9e36 (
    .a(al_615e209b[5]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[5]),
    .d(al_48cbf9af),
    .e(al_e890342d[5]),
    .o(al_ba2f1510[5]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_3cc211b7 (
    .a(al_615e209b[6]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[6]),
    .d(al_48cbf9af),
    .e(al_e890342d[6]),
    .o(al_ba2f1510[6]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_f49f1ee8 (
    .a(al_615e209b[7]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[7]),
    .d(al_48cbf9af),
    .e(al_e890342d[7]),
    .o(al_ba2f1510[7]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_a7bf881e (
    .a(al_615e209b[8]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[8]),
    .d(al_48cbf9af),
    .e(al_e890342d[8]),
    .o(al_ba2f1510[8]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(C)*~(D)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*~(D)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*C*D+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*C*D)"),
    .INIT(32'hf0eef022))
    al_d17e172a (
    .a(al_615e209b[9]),
    .b(al_d6af4c70[17]),
    .c(al_e8eb449b[9]),
    .d(al_48cbf9af),
    .e(al_e890342d[9]),
    .o(al_ba2f1510[9]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_75abaab7 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[14]),
    .c(al_f178cf22[15]),
    .o(al_64522de4));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'h5f5c5350))
    al_83306c16 (
    .a(al_489ab129),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[4]),
    .e(al_f178cf22[5]),
    .o(al_c18c443d));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'h5f5c5350))
    al_f293abe3 (
    .a(al_6bd097c8),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[8]),
    .e(al_f178cf22[9]),
    .o(al_63f07c7f));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_e30c6cb0 (
    .a(al_f120ad54),
    .b(al_63f07c7f),
    .c(al_b029b709[2]),
    .o(al_e54f5937));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7e233a00 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[0]),
    .c(al_f178cf22[1]),
    .o(al_267693c3));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*~(A)*~(E)+~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*A*~(E)+~(~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))*A*E+~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*A*E)"),
    .INIT(32'haaaa33f0))
    al_b885919f (
    .a(al_c18c443d),
    .b(al_d32b8d83),
    .c(al_267693c3),
    .d(al_b029b709[1]),
    .e(al_b029b709[2]),
    .o(al_f2ea1b91));
  AL_MAP_LUT5 #(
    .EQN("~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*~(C)*~(E)+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*~(E)+~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))*C*E+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*E)"),
    .INIT(32'h0f0f55cc))
    al_e2f60b7e (
    .a(al_e54f5937),
    .b(al_f2ea1b91),
    .c(al_c03651db),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_b0aa8206[0]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_71a13c13 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[10]),
    .c(al_f178cf22[11]),
    .o(al_6bd097c8));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'h5f5c5350))
    al_2490363a (
    .a(al_64522de4),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[12]),
    .e(al_f178cf22[13]),
    .o(al_f120ad54));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_c7d16c7d (
    .a(al_b029b709[0]),
    .b(al_f178cf22[6]),
    .c(al_f178cf22[7]),
    .o(al_489ab129));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_49672dc1 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[2]),
    .c(al_f178cf22[3]),
    .o(al_d32b8d83));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bc7ed73 (
    .a(al_b5005b7),
    .b(al_cd305354),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[10]));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))*~(C)+~E*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*~(C)+~(~E)*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C+~E*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C)"),
    .INIT(32'h5fcf50c0))
    al_3015d666 (
    .a(al_4ab15cc0),
    .b(al_c41ea483),
    .c(al_cd305354),
    .d(al_b029b709[2]),
    .e(al_f178cf22[17]),
    .o(al_b0aa8206[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_c2a9e609 (
    .a(al_40edf471),
    .b(al_cd305354),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[12]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A)*~((~C*B))+D*A*~((~C*B))+~(D)*A*(~C*B)+D*A*(~C*B))"),
    .INIT(16'hfb08))
    al_67302a88 (
    .a(al_14d0775),
    .b(al_cd305354),
    .c(al_b029b709[2]),
    .d(al_f178cf22[17]),
    .o(al_b0aa8206[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_bb859c52 (
    .a(al_e0531380),
    .b(al_cd305354),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_afb9f081 (
    .a(al_3c344131),
    .b(al_cd305354),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[15]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_5e6fcf5d (
    .a(al_b029b709[0]),
    .b(al_b029b709[1]),
    .o(al_5a076585));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_c42e927b (
    .a(al_b029b709[2]),
    .b(al_b029b709[3]),
    .o(al_1ce14aac));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    al_ea39cbb9 (
    .a(al_5a076585),
    .b(al_f178cf22[16]),
    .c(al_f178cf22[17]),
    .o(al_854c573f));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    al_d196e862 (
    .a(al_854c573f),
    .b(al_1ce14aac),
    .c(al_f178cf22[17]),
    .o(al_c03651db));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    al_4727fdde (
    .a(al_c03651db),
    .b(al_b029b709[4]),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[16]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_d94f124 (
    .a(al_14d0775),
    .b(al_923aa1f3),
    .c(al_b029b709[2]),
    .o(al_e841d7a8));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_5f897aaa (
    .a(al_88f2b0ea),
    .b(al_b029b709[2]),
    .o(al_e08923c5));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    al_7c9de39 (
    .a(al_c04f33dd),
    .b(al_b029b709[0]),
    .c(al_f178cf22[1]),
    .d(al_f178cf22[2]),
    .o(al_45f63f66));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    al_4db5effd (
    .a(al_45f63f66),
    .b(al_abf6101b),
    .c(al_cd305354),
    .d(al_86baf6c6),
    .o(al_5072ec3a));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~B)*~(D*A))"),
    .INIT(32'h000045cf))
    al_546bc401 (
    .a(al_e841d7a8),
    .b(al_e08923c5),
    .c(al_5072ec3a),
    .d(al_73eda6f6),
    .e(al_747e69b3),
    .o(al_b0aa8206[1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_af84b328 (
    .a(al_ab37028c),
    .b(al_185cfc7b),
    .c(al_b029b709[2]),
    .o(al_b5005b7));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_fc126d11 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[4]),
    .c(al_f178cf22[5]),
    .o(al_895351d0));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(E)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(E)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*E+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*E)"),
    .INIT(32'haaaa330f))
    al_d57823bd (
    .a(al_2b296468),
    .b(al_895351d0),
    .c(al_d32b8d83),
    .d(al_b029b709[1]),
    .e(al_b029b709[2]),
    .o(al_4c309c76));
  AL_MAP_LUT5 #(
    .EQN("(~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)*~(E)*~(D)+~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)*E*~(D)+~(~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))*E*D+~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)*E*D)"),
    .INIT(32'hff5c005c))
    al_e65e538f (
    .a(al_b5005b7),
    .b(al_4c309c76),
    .c(al_b029b709[3]),
    .d(al_b029b709[4]),
    .e(al_f178cf22[17]),
    .o(al_b0aa8206[2]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'h2e))
    al_cc75f0aa (
    .a(al_8a394456),
    .b(al_b029b709[1]),
    .c(al_f178cf22[17]),
    .o(al_4ab15cc0));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*~B))"),
    .INIT(16'h4050))
    al_44330a2c (
    .a(al_75f92221),
    .b(al_abf6101b),
    .c(al_cd305354),
    .d(al_c04f33dd),
    .o(al_60b812b4));
  AL_MAP_LUT5 #(
    .EQN("(~D*~A*~(B*~(E*C)))"),
    .INIT(32'h00510011))
    al_c7da231e (
    .a(al_a26df073),
    .b(al_60b812b4),
    .c(al_9ea7dc42),
    .d(al_747e69b3),
    .e(al_b029b709[2]),
    .o(al_b0aa8206[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_89888e49 (
    .a(al_b029b709[1]),
    .b(al_b029b709[2]),
    .o(al_86baf6c6));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_e83305b5 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[3]),
    .c(al_f178cf22[4]),
    .o(al_abf6101b));
  AL_MAP_LUT4 #(
    .EQN("(C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'ha030))
    al_262c72a9 (
    .a(al_4ab15cc0),
    .b(al_c41ea483),
    .c(al_73eda6f6),
    .d(al_b029b709[2]),
    .o(al_a26df073));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    al_2c12f4b6 (
    .a(al_86baf6c6),
    .b(al_b029b709[0]),
    .c(al_f178cf22[5]),
    .d(al_f178cf22[6]),
    .o(al_75f92221));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    al_c7f0c92c (
    .a(al_f120ad54),
    .b(al_854c573f),
    .c(al_b029b709[2]),
    .o(al_40edf471));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d0e9fde0 (
    .a(al_c18c443d),
    .b(al_63f07c7f),
    .c(al_b029b709[2]),
    .o(al_e7e648ec));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_9a37c04b (
    .a(al_e7e648ec),
    .b(al_40edf471),
    .c(al_b029b709[3]),
    .d(al_b029b709[4]),
    .e(al_f178cf22[17]),
    .o(al_b0aa8206[4]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'h5f5c5350))
    al_4c4617be (
    .a(al_8a394456),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[13]),
    .e(al_f178cf22[14]),
    .o(al_14d0775));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    al_9e53c93f (
    .a(al_9047c71),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[11]),
    .e(al_f178cf22[12]),
    .o(al_923aa1f3));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(A)*~(C)+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*~(C)+~(~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*A*C+~(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*A*C)"),
    .INIT(32'h5f5c5350))
    al_964ac45b (
    .a(al_9800fd32),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[5]),
    .e(al_f178cf22[6]),
    .o(al_88f2b0ea));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h10d0))
    al_5fbfa66f (
    .a(al_14d0775),
    .b(al_b029b709[2]),
    .c(al_b029b709[3]),
    .d(al_f178cf22[17]),
    .o(al_87b4efd6));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    al_500b7 (
    .a(al_923aa1f3),
    .b(al_88f2b0ea),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_1f3b4767));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    al_67c8e95d (
    .a(al_1f3b4767),
    .b(al_87b4efd6),
    .c(al_b029b709[4]),
    .d(al_f178cf22[17]),
    .o(al_b0aa8206[5]));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    al_6dd73d6 (
    .a(al_64522de4),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[16]),
    .e(al_f178cf22[17]),
    .o(al_ab37028c));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    al_e5d48500 (
    .a(al_6bd097c8),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[12]),
    .e(al_f178cf22[13]),
    .o(al_185cfc7b));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    al_7c0e128e (
    .a(al_ab37028c),
    .b(al_b029b709[2]),
    .c(al_f178cf22[17]),
    .o(al_e0531380));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    al_c35e0730 (
    .a(al_489ab129),
    .b(al_b029b709[0]),
    .c(al_b029b709[1]),
    .d(al_f178cf22[8]),
    .e(al_f178cf22[9]),
    .o(al_2b296468));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    al_6f2fbb85 (
    .a(al_185cfc7b),
    .b(al_2b296468),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_af16dfa7));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(C*~B))*~(E)*~(D)+(~A*~(C*~B))*E*~(D)+~((~A*~(C*~B)))*E*D+(~A*~(C*~B))*E*D)"),
    .INIT(32'hff450045))
    al_86a0881d (
    .a(al_af16dfa7),
    .b(al_e0531380),
    .c(al_b029b709[3]),
    .d(al_b029b709[4]),
    .e(al_f178cf22[17]),
    .o(al_b0aa8206[6]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_57c47d79 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[15]),
    .c(al_f178cf22[16]),
    .o(al_8a394456));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_a7c0acce (
    .a(al_9047c71),
    .b(al_9800fd32),
    .c(al_b029b709[1]),
    .o(al_9ea7dc42));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a45b5890 (
    .a(al_9ea7dc42),
    .b(al_c41ea483),
    .c(al_b029b709[2]),
    .o(al_879333c8));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*~(E)*~(D)+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*~(D)+~((A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))*E*D+(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)*E*D)"),
    .INIT(32'hffca00ca))
    al_6aecfd27 (
    .a(al_879333c8),
    .b(al_3c344131),
    .c(al_b029b709[3]),
    .d(al_b029b709[4]),
    .e(al_f178cf22[17]),
    .o(al_b0aa8206[7]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_da186c54 (
    .a(al_b029b709[0]),
    .b(al_f178cf22[9]),
    .c(al_f178cf22[10]),
    .o(al_9047c71));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    al_fc5ecb93 (
    .a(al_f178cf22[14]),
    .b(al_f178cf22[13]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_1259ba86));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_3a6c9a75 (
    .a(al_f178cf22[11]),
    .b(al_f178cf22[12]),
    .c(al_1259ba86),
    .d(al_b029b709[1]),
    .o(al_c41ea483));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_3953e9ef (
    .a(al_8a394456),
    .b(al_c04f33dd),
    .c(al_f178cf22[17]),
    .o(al_3c344131));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    al_75c7e8ff (
    .a(al_b029b709[0]),
    .b(al_f178cf22[7]),
    .c(al_f178cf22[8]),
    .o(al_9800fd32));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_3f463ee5 (
    .a(al_b029b709[3]),
    .b(al_b029b709[4]),
    .o(al_73eda6f6));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_c7a21ab1 (
    .a(al_b029b709[4]),
    .b(al_f178cf22[17]),
    .o(al_747e69b3));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E)"),
    .INIT(32'h00f8fcf8))
    al_529237a1 (
    .a(al_854c573f),
    .b(al_73eda6f6),
    .c(al_747e69b3),
    .d(al_b029b709[2]),
    .e(al_f178cf22[17]),
    .o(al_51f316f6));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    al_1e979d92 (
    .a(al_e54f5937),
    .b(al_51f316f6),
    .c(al_cd305354),
    .o(al_b0aa8206[8]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_bf0b8ab (
    .a(al_e841d7a8),
    .b(al_cd305354),
    .c(al_f178cf22[17]),
    .o(al_b0aa8206[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_17f09c3c (
    .a(al_5f6ba172),
    .b(xin[0]),
    .c(yin[0]),
    .o(al_8b1ee5d9[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4c8e5fdd (
    .a(al_5f6ba172),
    .b(xin[10]),
    .c(yin[10]),
    .o(al_8b1ee5d9[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_12078e2f (
    .a(al_5f6ba172),
    .b(xin[11]),
    .c(yin[11]),
    .o(al_8b1ee5d9[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d5590079 (
    .a(al_5f6ba172),
    .b(xin[12]),
    .c(yin[12]),
    .o(al_8b1ee5d9[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_7fd7472e (
    .a(al_5f6ba172),
    .b(xin[13]),
    .c(yin[13]),
    .o(al_8b1ee5d9[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_22f8cd3e (
    .a(al_5f6ba172),
    .b(xin[14]),
    .c(yin[14]),
    .o(al_8b1ee5d9[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f5fe3baf (
    .a(al_5f6ba172),
    .b(xin[15]),
    .c(yin[15]),
    .o(al_8b1ee5d9[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f3ebe195 (
    .a(al_5f6ba172),
    .b(xin[16]),
    .c(yin[16]),
    .o(al_8b1ee5d9[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_66c388a6 (
    .a(al_5f6ba172),
    .b(xin[1]),
    .c(yin[1]),
    .o(al_8b1ee5d9[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a6a60456 (
    .a(al_5f6ba172),
    .b(xin[2]),
    .c(yin[2]),
    .o(al_8b1ee5d9[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_6e9130ae (
    .a(al_5f6ba172),
    .b(xin[3]),
    .c(yin[3]),
    .o(al_8b1ee5d9[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_bb990db6 (
    .a(xin[17]),
    .b(yin[17]),
    .o(al_5f6ba172));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_1a017fe (
    .a(al_5f6ba172),
    .b(xin[4]),
    .c(yin[4]),
    .o(al_8b1ee5d9[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_fcdeeda7 (
    .a(al_5f6ba172),
    .b(xin[5]),
    .c(yin[5]),
    .o(al_8b1ee5d9[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4dbeb136 (
    .a(al_5f6ba172),
    .b(xin[6]),
    .c(yin[6]),
    .o(al_8b1ee5d9[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b62a2eec (
    .a(al_5f6ba172),
    .b(xin[7]),
    .c(yin[7]),
    .o(al_8b1ee5d9[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4c02872e (
    .a(al_5f6ba172),
    .b(xin[8]),
    .c(yin[8]),
    .o(al_8b1ee5d9[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_2b8706cf (
    .a(al_5f6ba172),
    .b(xin[9]),
    .c(yin[9]),
    .o(al_8b1ee5d9[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_61996160 (
    .a(al_83a98034),
    .b(al_f774eaf9[0]),
    .c(al_655add9[0]),
    .o(al_7b6549fa[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_8a0ea400 (
    .a(al_83a98034),
    .b(al_54f6e7c3[10]),
    .c(al_f774eaf9[10]),
    .o(al_7b6549fa[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_97085dca (
    .a(al_83a98034),
    .b(al_54f6e7c3[11]),
    .c(al_f774eaf9[11]),
    .o(al_7b6549fa[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c08a7b95 (
    .a(al_83a98034),
    .b(al_54f6e7c3[12]),
    .c(al_f774eaf9[12]),
    .o(al_7b6549fa[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_408266ea (
    .a(al_83a98034),
    .b(al_54f6e7c3[13]),
    .c(al_f774eaf9[13]),
    .o(al_7b6549fa[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_c8be92ee (
    .a(al_83a98034),
    .b(al_54f6e7c3[14]),
    .c(al_f774eaf9[14]),
    .o(al_7b6549fa[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3b15e97e (
    .a(al_83a98034),
    .b(al_54f6e7c3[15]),
    .c(al_f774eaf9[15]),
    .o(al_7b6549fa[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_26823686 (
    .a(al_83a98034),
    .b(al_54f6e7c3[16]),
    .c(al_f774eaf9[16]),
    .o(al_7b6549fa[16]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    al_a2a1a5e (
    .a(al_54f6e7c3[17]),
    .b(al_f774eaf9[17]),
    .c(al_655add9[17]),
    .o(al_7b6549fa[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_43db0c91 (
    .a(al_83a98034),
    .b(al_54f6e7c3[1]),
    .c(al_f774eaf9[1]),
    .o(al_7b6549fa[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_633c6224 (
    .a(al_83a98034),
    .b(al_54f6e7c3[2]),
    .c(al_f774eaf9[2]),
    .o(al_7b6549fa[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d36f09f0 (
    .a(al_83a98034),
    .b(al_54f6e7c3[3]),
    .c(al_f774eaf9[3]),
    .o(al_7b6549fa[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_bae032d3 (
    .a(al_83a98034),
    .b(al_54f6e7c3[4]),
    .c(al_f774eaf9[4]),
    .o(al_7b6549fa[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_96d8146c (
    .a(al_83a98034),
    .b(al_54f6e7c3[5]),
    .c(al_f774eaf9[5]),
    .o(al_7b6549fa[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3ebfa08c (
    .a(al_83a98034),
    .b(al_54f6e7c3[6]),
    .c(al_f774eaf9[6]),
    .o(al_7b6549fa[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_51faf1d5 (
    .a(al_83a98034),
    .b(al_54f6e7c3[7]),
    .c(al_f774eaf9[7]),
    .o(al_7b6549fa[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_aa1ca45b (
    .a(al_83a98034),
    .b(al_54f6e7c3[8]),
    .c(al_f774eaf9[8]),
    .o(al_7b6549fa[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_281d9e01 (
    .a(al_83a98034),
    .b(al_54f6e7c3[9]),
    .c(al_f774eaf9[9]),
    .o(al_7b6549fa[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_da1d08f (
    .a(al_9a3f7017[0]),
    .b(al_12c226aa[0]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[0]),
    .o(al_a89eb1ca[0]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_e71a1331 (
    .a(al_9a3f7017[10]),
    .b(al_12c226aa[10]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[10]),
    .o(al_a89eb1ca[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_b00fbc02 (
    .a(al_9a3f7017[11]),
    .b(al_12c226aa[11]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[11]),
    .o(al_a89eb1ca[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_e03e8b2 (
    .a(al_9a3f7017[12]),
    .b(al_12c226aa[12]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[12]),
    .o(al_a89eb1ca[12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_21ae4b3e (
    .a(al_9a3f7017[13]),
    .b(al_12c226aa[13]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[13]),
    .o(al_a89eb1ca[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_a733c5a6 (
    .a(al_9a3f7017[14]),
    .b(al_12c226aa[14]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[14]),
    .o(al_a89eb1ca[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_c45a8ef0 (
    .a(al_9a3f7017[15]),
    .b(al_12c226aa[15]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[15]),
    .o(al_a89eb1ca[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_1db5572f (
    .a(al_9a3f7017[16]),
    .b(al_12c226aa[16]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[16]),
    .o(al_a89eb1ca[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_d723e4c4 (
    .a(al_9a3f7017[17]),
    .b(al_12c226aa[17]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[17]),
    .o(al_a89eb1ca[17]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_64ae39a3 (
    .a(al_9a3f7017[1]),
    .b(al_12c226aa[1]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[1]),
    .o(al_a89eb1ca[1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_1193e73c (
    .a(al_9a3f7017[2]),
    .b(al_12c226aa[2]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[2]),
    .o(al_a89eb1ca[2]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_2691f80d (
    .a(al_9a3f7017[3]),
    .b(al_12c226aa[3]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[3]),
    .o(al_a89eb1ca[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_42d825ad (
    .a(al_9a3f7017[4]),
    .b(al_12c226aa[4]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[4]),
    .o(al_a89eb1ca[4]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_ae92dfee (
    .a(al_9a3f7017[5]),
    .b(al_12c226aa[5]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[5]),
    .o(al_a89eb1ca[5]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_8b959a59 (
    .a(al_9a3f7017[6]),
    .b(al_12c226aa[6]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[6]),
    .o(al_a89eb1ca[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_96aaf6c (
    .a(al_9a3f7017[7]),
    .b(al_12c226aa[7]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[7]),
    .o(al_a89eb1ca[7]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_5b3b424d (
    .a(al_9a3f7017[8]),
    .b(al_12c226aa[8]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[8]),
    .o(al_a89eb1ca[8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(B)*~(D)+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*~(D)+~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*B*D+(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*B*D)"),
    .INIT(32'hccafcca0))
    al_6a1c2d53 (
    .a(al_9a3f7017[9]),
    .b(al_12c226aa[9]),
    .c(al_d6af4c70[17]),
    .d(al_48cbf9af),
    .e(al_deeec3ed[9]),
    .o(al_a89eb1ca[9]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_ba6dee4a (
    .a(al_d6af4c70[10]),
    .b(al_d6af4c70[11]),
    .c(al_b029b709[0]),
    .o(al_248f265c));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'h5555f0cc))
    al_4de182d (
    .a(al_1de057dc),
    .b(al_d6af4c70[4]),
    .c(al_d6af4c70[5]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_dee61509));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'h5555f0cc))
    al_b94e84ca (
    .a(al_248f265c),
    .b(al_d6af4c70[8]),
    .c(al_d6af4c70[9]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_ce078ee));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_b5e81755 (
    .a(al_2b0d498c),
    .b(al_ce078ee),
    .c(al_b029b709[2]),
    .o(al_6652589d));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    al_eff1cf2b (
    .a(al_329701d8),
    .b(al_d6af4c70[17]),
    .c(al_b029b709[3]),
    .d(al_b029b709[4]),
    .o(al_9aa2c63b));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9258a21d (
    .a(al_d6af4c70[0]),
    .b(al_d6af4c70[1]),
    .c(al_b029b709[0]),
    .o(al_44f78eb0));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*~(A)*~(E)+~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*A*~(E)+~(~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))*A*E+~(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D)*A*E)"),
    .INIT(32'haaaa33f0))
    al_a7e5efb (
    .a(al_dee61509),
    .b(al_399025e4),
    .c(al_44f78eb0),
    .d(al_b029b709[1]),
    .e(al_b029b709[2]),
    .o(al_b494668c));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)))"),
    .INIT(32'hf0f0f5fc))
    al_d240ef70 (
    .a(al_6652589d),
    .b(al_b494668c),
    .c(al_9aa2c63b),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_9addee19[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    al_f048e819 (
    .a(al_d6af4c70[14]),
    .b(al_d6af4c70[15]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_efe81361));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_203a84a5 (
    .a(al_d6af4c70[12]),
    .b(al_d6af4c70[13]),
    .c(al_efe81361),
    .d(al_b029b709[1]),
    .o(al_2b0d498c));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_93633271 (
    .a(al_d6af4c70[6]),
    .b(al_d6af4c70[7]),
    .c(al_b029b709[0]),
    .o(al_1de057dc));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_deadbbfd (
    .a(al_d6af4c70[2]),
    .b(al_d6af4c70[3]),
    .c(al_b029b709[0]),
    .o(al_399025e4));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    al_4adda60e (
    .a(al_967be913),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .o(al_9addee19[10]));
  AL_MAP_LUT5 #(
    .EQN("(D*~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*~(C)+D*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)+~(D)*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C+D*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C)"),
    .INIT(32'hcfc0afa0))
    al_dc097297 (
    .a(al_2853bf2a),
    .b(al_ce27e68f),
    .c(al_cd305354),
    .d(al_d6af4c70[17]),
    .e(al_b029b709[2]),
    .o(al_9addee19[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_455a96f7 (
    .a(al_5f96adf7),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .o(al_9addee19[12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A)*~((~D*B))+C*A*~((~D*B))+~(C)*A*(~D*B)+C*A*(~D*B))"),
    .INIT(16'hf0b8))
    al_a1dbe7c5 (
    .a(al_c29dd627),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[2]),
    .o(al_9addee19[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_2444681 (
    .a(al_31cf9bca),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .o(al_9addee19[14]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A)*~((~D*B))+C*A*~((~D*B))+~(C)*A*(~D*B)+C*A*(~D*B))"),
    .INIT(16'hf0b8))
    al_7e099f62 (
    .a(al_ce27e68f),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[2]),
    .o(al_9addee19[15]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((~D*A))+C*B*~((~D*A))+~(C)*B*(~D*A)+C*B*(~D*A))"),
    .INIT(16'hf0d8))
    al_3d749278 (
    .a(al_5a076585),
    .b(al_d6af4c70[16]),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[2]),
    .o(al_329701d8));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    al_b78fcc0d (
    .a(al_329701d8),
    .b(al_cd305354),
    .c(al_d6af4c70[17]),
    .o(al_9addee19[16]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h5300))
    al_41c1c8b0 (
    .a(al_c29dd627),
    .b(al_d92048f7),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_fb209166));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    al_37338b62 (
    .a(al_d6af4c70[1]),
    .b(al_d6af4c70[2]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_b77cbcd0));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    al_a5edab96 (
    .a(al_d6af4c70[3]),
    .b(al_d6af4c70[4]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_6075e6a9));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .INIT(32'h000055fc))
    al_43e32840 (
    .a(al_9ca1c07c),
    .b(al_b77cbcd0),
    .c(al_6075e6a9),
    .d(al_b029b709[2]),
    .e(al_b029b709[3]),
    .o(al_492fb484));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(C)*~(D)+(~B*~A)*C*~(D)+~((~B*~A))*C*D+(~B*~A)*C*D)"),
    .INIT(16'hf011))
    al_aced97fd (
    .a(al_fb209166),
    .b(al_492fb484),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[4]),
    .o(al_9addee19[1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_1a8c54ef (
    .a(al_85347eda),
    .b(al_96795d02),
    .c(al_b029b709[2]),
    .o(al_967be913));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_db741694 (
    .a(al_d6af4c70[4]),
    .b(al_d6af4c70[5]),
    .c(al_b029b709[0]),
    .o(al_dce5c03c));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_609615d8 (
    .a(al_dce5c03c),
    .b(al_399025e4),
    .c(al_b029b709[1]),
    .d(al_b029b709[2]),
    .o(al_48b19352));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    al_7fd179c1 (
    .a(al_598dbbb7),
    .b(al_1de057dc),
    .c(al_48b19352),
    .d(al_b029b709[2]),
    .o(al_6af624ab));
  AL_MAP_LUT5 #(
    .EQN("(~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*~(C)*~(E)+~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*~(E)+~(~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))*C*E+~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*E)"),
    .INIT(32'hf0f055cc))
    al_e05f7e84 (
    .a(al_967be913),
    .b(al_6af624ab),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_9addee19[2]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_15b42a43 (
    .a(al_d6af4c70[5]),
    .b(al_d6af4c70[6]),
    .c(al_b029b709[0]),
    .o(al_2013c010));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(A)*~(E)+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*~(E)+~(~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*A*E+~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*A*E)"),
    .INIT(32'haaaa0f33))
    al_39cfa3ec (
    .a(al_2013c010),
    .b(al_d6af4c70[3]),
    .c(al_d6af4c70[4]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_22d6ddd));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~B)*~(~C*~A))"),
    .INIT(16'hfac8))
    al_93633882 (
    .a(al_f42f533c),
    .b(al_22d6ddd),
    .c(al_1ce14aac),
    .d(al_b029b709[2]),
    .o(al_b5596380));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    al_ce88be1c (
    .a(al_2853bf2a),
    .b(al_ce27e68f),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_65737be6));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(C)*~(D)+(~B*~A)*C*~(D)+~((~B*~A))*C*D+(~B*~A)*C*D)"),
    .INIT(16'hf011))
    al_fbbe762a (
    .a(al_b5596380),
    .b(al_65737be6),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[4]),
    .o(al_9addee19[3]));
  AL_MAP_LUT5 #(
    .EQN("(A*~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*~(E)+A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(E)+~(A)*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*E+A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*E)"),
    .INIT(32'hf3c0aaaa))
    al_cff1964b (
    .a(al_2b0d498c),
    .b(al_5a076585),
    .c(al_d6af4c70[16]),
    .d(al_d6af4c70[17]),
    .e(al_b029b709[2]),
    .o(al_5f96adf7));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2f5ec807 (
    .a(al_dee61509),
    .b(al_ce078ee),
    .c(al_b029b709[2]),
    .o(al_1883443));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*~(C)*~(E)+(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*C*~(E)+~((A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))*C*E+(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*C*E)"),
    .INIT(32'hf0f0ccaa))
    al_11d70bed (
    .a(al_1883443),
    .b(al_5f96adf7),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_9addee19[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    al_bfd658fd (
    .a(al_d6af4c70[15]),
    .b(al_d6af4c70[16]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_1fb8f7d6));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(C)*~(D)+(~B*~A)*C*~(D)+~((~B*~A))*C*D+(~B*~A)*C*D)"),
    .INIT(16'hf011))
    al_b211f57 (
    .a(al_6d3f1d3d),
    .b(al_137b074e),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[4]),
    .o(al_9addee19[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_45aae0af (
    .a(al_d6af4c70[13]),
    .b(al_d6af4c70[14]),
    .c(al_1fb8f7d6),
    .d(al_b029b709[1]),
    .o(al_c29dd627));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E)"),
    .INIT(32'hf0cc5555))
    al_7ecb0aca (
    .a(al_72ad6500),
    .b(al_d6af4c70[11]),
    .c(al_d6af4c70[12]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_d92048f7));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E)"),
    .INIT(32'hf0cc5555))
    al_404601e9 (
    .a(al_2013c010),
    .b(al_d6af4c70[7]),
    .c(al_d6af4c70[8]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_9ca1c07c));
  AL_MAP_LUT4 #(
    .EQN("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h3500))
    al_9d1902ea (
    .a(al_c29dd627),
    .b(al_d6af4c70[17]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_137b074e));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h0053))
    al_45ecf308 (
    .a(al_d92048f7),
    .b(al_9ca1c07c),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_6d3f1d3d));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    al_7ba702e6 (
    .a(al_d6af4c70[16]),
    .b(al_d6af4c70[17]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_6c78c52c));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(D*~B))*~(C)*~(E)+(~A*~(D*~B))*C*~(E)+~((~A*~(D*~B)))*C*E+(~A*~(D*~B))*C*E)"),
    .INIT(32'hf0f04455))
    al_c67f4861 (
    .a(al_a2275c94),
    .b(al_31cf9bca),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_9addee19[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_77da14d3 (
    .a(al_d6af4c70[14]),
    .b(al_d6af4c70[15]),
    .c(al_6c78c52c),
    .d(al_b029b709[1]),
    .o(al_85347eda));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))*~(E)+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*~(E)+~(~A)*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E+~A*(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)*E)"),
    .INIT(32'hf0cc5555))
    al_a669e9df (
    .a(al_248f265c),
    .b(al_d6af4c70[12]),
    .c(al_d6af4c70[13]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_96795d02));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ee717165 (
    .a(al_85347eda),
    .b(al_d6af4c70[17]),
    .c(al_b029b709[2]),
    .o(al_31cf9bca));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_d32f15fc (
    .a(al_d6af4c70[8]),
    .b(al_d6af4c70[9]),
    .c(al_b029b709[0]),
    .o(al_598dbbb7));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    al_a3f5b53b (
    .a(al_598dbbb7),
    .b(al_1de057dc),
    .c(al_b029b709[1]),
    .o(al_4772cc8e));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'h0035))
    al_354325d6 (
    .a(al_4772cc8e),
    .b(al_96795d02),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_a2275c94));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_62e44beb (
    .a(al_d6af4c70[9]),
    .b(al_d6af4c70[10]),
    .c(al_b029b709[0]),
    .o(al_72ad6500));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    al_a04111f2 (
    .a(al_72ad6500),
    .b(al_80739918),
    .c(al_b029b709[1]),
    .d(al_b029b709[3]),
    .o(al_f42f533c));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_b4f3b175 (
    .a(al_2853bf2a),
    .b(al_b029b709[3]),
    .o(al_853b0020));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)*~(D)*~(E)+~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)*D*~(E)+~(~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B))*D*E+~(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)*D*E)"),
    .INIT(32'hff002e2e))
    al_295a7277 (
    .a(al_853b0020),
    .b(al_67d43207),
    .c(al_f42f533c),
    .d(al_d6af4c70[17]),
    .e(al_b029b709[4]),
    .o(al_9addee19[7]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*~(C)*~(E)+(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*C*~(E)+~((A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))*C*E+(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)*C*E)"),
    .INIT(32'hf0f0ccaa))
    al_c66dcfd7 (
    .a(al_d6af4c70[15]),
    .b(al_d6af4c70[16]),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[0]),
    .e(al_b029b709[1]),
    .o(al_ce27e68f));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    al_29b26a3a (
    .a(al_d6af4c70[13]),
    .b(al_d6af4c70[14]),
    .c(al_b029b709[0]),
    .d(al_b029b709[1]),
    .o(al_b2a8a0cc));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    al_5b936a11 (
    .a(al_d6af4c70[11]),
    .b(al_d6af4c70[12]),
    .c(al_b2a8a0cc),
    .d(al_b029b709[1]),
    .o(al_2853bf2a));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    al_922b5dcc (
    .a(al_d6af4c70[7]),
    .b(al_d6af4c70[8]),
    .c(al_b029b709[0]),
    .o(al_80739918));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    al_9fb1eef8 (
    .a(al_ce27e68f),
    .b(al_d6af4c70[17]),
    .c(al_b029b709[2]),
    .d(al_b029b709[3]),
    .o(al_67d43207));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D)*~(C)*~(E)+(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D)*C*~(E)+~((~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))*C*E+(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D)*C*E)"),
    .INIT(32'hf0f0cc55))
    al_9d867aea (
    .a(al_6652589d),
    .b(al_329701d8),
    .c(al_d6af4c70[17]),
    .d(al_b029b709[3]),
    .e(al_b029b709[4]),
    .o(al_9addee19[8]));
  AL_MAP_LUT5 #(
    .EQN("(D*~((B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E))*~(C)+D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)*~(C)+~(D)*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)*C+D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)*C)"),
    .INIT(32'hafa0cfc0))
    al_936d0d05 (
    .a(al_c29dd627),
    .b(al_d92048f7),
    .c(al_cd305354),
    .d(al_d6af4c70[17]),
    .e(al_b029b709[2]),
    .o(al_9addee19[9]));

endmodule 

