module calculate (
    input wire clk,
    input wire rstn,
    input wire [16: 0] real1,
    input wire [16: 0] image1,

    output wire [15: 0] r_out,
    output wire [15: 0] z_out
);

//assign r_out = () / ();
//assign z_out = 

endmodule